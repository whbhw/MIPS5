`define NOP_INST        32'h0000_0020
`define NOP_CTRL        16'b010_0000110100000
`define NOP_MEM_CTRL    6'b000010
`define NOP_WB_CTRL     4'b0010

`define DEFAULT_PC      32'h_00400000
`define DEFAULT_PC_4    32'h_00400004