`define INST_NOP 32'h0000_0020
`define DEFAULT_PC 32'h_00400000
`define DEFAULT_PC_4 32'h_00400004