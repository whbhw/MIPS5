module EXTEND (
    output  wire    [31:0]  extend_out  ,
    input   wire    [15:0]  extend_in   ,
    input   wire            signext     
);

endmodule